library verilog;
use verilog.vl_types.all;
entity CNT_of_rattle_vlg_vec_tst is
end CNT_of_rattle_vlg_vec_tst;
