library verilog;
use verilog.vl_types.all;
entity SchematicStatus_vlg_vec_tst is
end SchematicStatus_vlg_vec_tst;
