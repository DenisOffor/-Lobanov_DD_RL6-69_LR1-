library verilog;
use verilog.vl_types.all;
entity Code_converter_vlg_vec_tst is
end Code_converter_vlg_vec_tst;
