library verilog;
use verilog.vl_types.all;
entity SyncCNT_vlg_vec_tst is
end SyncCNT_vlg_vec_tst;
